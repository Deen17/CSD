`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    
// Design Name: 
// Module Name:    loopback 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module loopback( switches, leds, rs232_tx, rs232_rx, reset, clk, col, row );

	// Top-level Inputs and Outputs
	// These connect directly to FPGA pins via the pin map
	//
	// Control - clk, rst, etc
	input			reset;			// Remember: ACTIVE LOW!!!
	input			clk;			// 100 MHz
	// GPIO
	input	[7:0]	switches;
	output	[7:0]	leds;
	// RS232 Lines
	input			rs232_rx;
	output			rs232_tx;
	
	//keypad
	output [3:0] col;
	input [3:0] row;
	
	// Wires and Register Declarations
	//
	// PicoBlaze Data Lines
	wire	[7:0]	pb_port_id;
	wire	[7:0]	pb_out_port;
	reg		[7:0]	pb_in_port;
	wire			pb_read_strobe;
	wire			pb_write_strobe;
	// PicoBlaze CPU Control Wires
	wire			pb_reset;
	wire			pb_interrupt;
	wire			pb_int_ack;
	
	// UART wires
	wire			write_to_uart;
	wire			uart_buffer_full;
	wire			uart_data_present;
	reg				read_from_uart;
	wire			uart_reset;
	// UART Data Lines
	// TX does not need a wire, as it is fed directly by pb_out_port
	wire	[7:0]	uart_rx_data;
	
	// LED wires
	wire write_to_leds;
	wire led_reset;
	

	// LED Driver and control logic
	//
	// LED driver expects ACTIVE-HIGH reset
	assign led_reset = reset;
	// LED driver instantiation
	led_driver_wrapper led_driver (
		.led_value(pb_out_port),
		.leds(leds),
		.write_to_leds(write_to_leds),
		.reset(led_reset),
		.clk(clk)
	);
	
	//keypad requires timer to shift col bits;
	wire [3:0] upc_out;

		up_counter upc(
			.clk(clk),
			.reset(reset),
			.out(upc_out)
		);
	assign col = upc_out;

	
	// UART and control logic
	//
	// UART expects ACTIVE-HIGH reset	
	assign uart_reset =  reset;
	// UART instantiation
	//
	// Within the UART Module (rs232_uart.v), make sure you fill in the
	// appropriate sections.
	rs232_uart UART (
		.tx_data_in(pb_out_port), // The UART only accepts data from PB, so we just tie the PB output to the UART input.
		.write_tx_data(write_to_uart), // Goes high when PB sends write strobe and PORT_ID is the UART write port number
		.tx_buffer_full(uart_buffer_full),
		.rx_data_out(uart_rx_data),
		.read_rx_data_ack(read_from_uart),
		.rx_data_present(uart_data_present),
		.rs232_tx(rs232_tx),
		.rs232_rx(rs232_rx),
		.reset(uart_reset),
		.clk(clk)
	);	
	
	// PicoBlaze and control logic
	//
	// PB expects ACTIVE-HIGH reset
	assign pb_reset = reset;
	// Disable interrupt by assigning 0 to interrupt
	assign pb_interrupt = 1'b0;
	// PB CPU instantiation
	//
	// Within the PicoBlaze Module (picoblaze.v), make sure you fill in the
	// appropriate sections.
	picoblaze CPU (
		.port_id(pb_port_id),
		.read_strobe(pb_read_strobe),
		.in_port(pb_in_port),
		.write_strobe(pb_write_strobe),
		.out_port(pb_out_port),
		.interrupt(pb_interrupt),
		.interrupt_ack(),
		.reset(pb_reset),
		.clk(clk)
	);	
	// PB I/O selection/routing
	//
	// Handle PicoBlaze Output Port Logic
	// Output Ports:
	// * leds_out : port 01
	// * uart_data_tx : port 03
	// * keys: port 06
	// 
	// These signals are effectively "write enable" lines for the UART and LED
	// Driver modules. They must be asserted when PB is outputting to the
	// corresponding port
	assign write_to_leds = pb_write_strobe & (pb_port_id == 8'h01);
	assign write_to_uart = pb_write_strobe & (pb_port_id == 8'h03 || pb_port_id == 8'h06);
	//
	// Handle PicoBlaze Input Port Logic
	// Input Ports:
	// * switches_in : port 00
	// * uart_data_rx : port 02
	// * uart_data_present : port 04 (1-bit, assigned to LSB)
	// * uart_buffer_full: port 05 (1-bit, assigned to LSB)
	//
	// This process block gets the value of the requested input port device
	// and passes it to PBs in_port. When PB is not requestng data from
	// a valid input port, set the input to static 0.
	reg [7:0] keyflag;
	always @(posedge clk or posedge pb_reset)
	begin
		if(pb_reset) begin
			pb_in_port <= 0;
			read_from_uart <= 0;
		end else begin
			// Set pb input port to appropriate value
			case(pb_port_id)
				8'h00: pb_in_port <= switches;
				8'h02: pb_in_port <= uart_rx_data; //waas uart_data_rx
				8'h04: pb_in_port <= {7'b0000000,uart_data_present};
				8'h05: pb_in_port <= {7'b0000000,uart_buffer_full};
				8'h06: pb_in_port <= keyflag;
				/*	begin
							if(!col[0] && !row[0]) begin
								pb_in_port <= 8'h01;
							end
							else if(!col[1] && !row[0]) begin
								pb_in_port <= 8'h02;
							end
							else if(!col[2] && !row[0]) begin
								pb_in_port <= 8'd03;
							end
							else if(!col[0] && !row[1]) begin
								pb_in_port <= 8'h04;
							end
							else if(!col[1] && !row[1]) begin
								pb_in_port <= 8'h05;
							end
							else begin
								pb_in_port <= 8'h0a;
							end
						end
*/				default: pb_in_port <= 8'h0a;
			endcase
			// Set up acknowledge/enable signals.
			//
			// Some modules, such as the UART, need confirmation that the data
			// has been read, since it needs to push it off the queue and make
			// the next byte available. This logic will set the 'read_from'
			// signal high for corresponding ports, as needed. Most input
			// ports will not need this.
			read_from_uart <= pb_read_strobe & (pb_port_id == 8'h04);
		end
	end
	
always @(posedge clk)
begin
	if(!col[0]&& !row[0])
		keyflag <= 8'h01;
	else if(!col[1]&& !row[0])
		keyflag <= 8'h02; 
	else if(!col[2]&& !row[0])
		keyflag <= 8'h03;
	else if(!col[0]&& !row[1])
		keyflag <= 8'h04;
	else if(!col[1]&& !row[1])
		keyflag <= 8'h05;
	else if(!col[2]&& !row[1])
		keyflag <= 8'h06;
	else if(!col[0]&& !row[2])
		keyflag <= 8'h07;
	else if(!col[1]&& !row[2])
		keyflag <= 8'h08;
	else if(!col[2]&& !row[2])
		keyflag <= 8'h09;
	else if(!col[0]&& !row[3])
		keyflag <= 8'h00;
	else if(!col[1]&& !row[3])
		keyflag <= 8'h0f;
	else if(!col[2]&& !row[3])
		keyflag <= 8'h0e;
	else if(!col[3]&& !row[0])
		keyflag <= 8'h0a;
	else if(!col[3]&& !row[1])
		keyflag <= 8'h0b;
	else if(!col[3]&& !row[2])
		keyflag <= 8'h0c;
	else if (!col[3]&&!row[3])
		keyflag <= 8'h0d;
	else keyflag <= 8'h00;
end

endmodule
